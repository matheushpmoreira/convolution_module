library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity convolution_module is

end convolution_module;

architecture arch of convolution_module is
begin
    
  
end arch;
